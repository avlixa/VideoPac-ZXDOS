-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d3",
     9 => x"98080b0b",
    10 => x"80d39c08",
    11 => x"0b0b80d3",
    12 => x"a0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d3a00c0b",
    16 => x"0b80d39c",
    17 => x"0c0b0b80",
    18 => x"d3980c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80c998",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d39870",
    57 => x"80ddd027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5196f1",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d3",
    65 => x"a80c9f0b",
    66 => x"80d3ac0c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d3ac08ff",
    70 => x"0580d3ac",
    71 => x"0c80d3ac",
    72 => x"088025e8",
    73 => x"3880d3a8",
    74 => x"08ff0580",
    75 => x"d3a80c80",
    76 => x"d3a80880",
    77 => x"25d03880",
    78 => x"0b80d3ac",
    79 => x"0c800b80",
    80 => x"d3a80c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d3a808",
   100 => x"25913882",
   101 => x"c82d80d3",
   102 => x"a808ff05",
   103 => x"80d3a80c",
   104 => x"838a0480",
   105 => x"d3a80880",
   106 => x"d3ac0853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d3a808",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d3ac0881",
   116 => x"0580d3ac",
   117 => x"0c80d3ac",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d3ac",
   121 => x"0c80d3a8",
   122 => x"08810580",
   123 => x"d3a80c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d3",
   128 => x"ac088105",
   129 => x"80d3ac0c",
   130 => x"80d3ac08",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d3ac",
   134 => x"0c80d3a8",
   135 => x"08810580",
   136 => x"d3a80c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d3b00cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"d3b00c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180d3",
   177 => x"b0088407",
   178 => x"80d3b00c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5485bc74",
   182 => x"258f3882",
   183 => x"0b0b0b80",
   184 => x"ce9c0c80",
   185 => x"d05385f3",
   186 => x"04810b0b",
   187 => x"0b80ce9c",
   188 => x"0cbc530b",
   189 => x"0b80ce9c",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0cfc0875",
   193 => x"7531ffb0",
   194 => x"05ff1371",
   195 => x"712cff94",
   196 => x"1a709f2a",
   197 => x"1170812c",
   198 => x"80d3b008",
   199 => x"52545153",
   200 => x"57535152",
   201 => x"5276802e",
   202 => x"85387081",
   203 => x"075170f6",
   204 => x"940c7209",
   205 => x"8105f680",
   206 => x"0c710981",
   207 => x"05f6840c",
   208 => x"0294050d",
   209 => x"0402f405",
   210 => x"0d745372",
   211 => x"70810554",
   212 => x"80f52d52",
   213 => x"71802e89",
   214 => x"38715183",
   215 => x"842d86cb",
   216 => x"04810b80",
   217 => x"d3980c02",
   218 => x"8c050d04",
   219 => x"02fc050d",
   220 => x"81808051",
   221 => x"c0115170",
   222 => x"fb380284",
   223 => x"050d0402",
   224 => x"fc050dec",
   225 => x"5183710c",
   226 => x"86ec2d82",
   227 => x"710c0284",
   228 => x"050d0486",
   229 => x"ec2d86ec",
   230 => x"2d86ec2d",
   231 => x"86ec2d86",
   232 => x"ec2d86ec",
   233 => x"2d86ec2d",
   234 => x"86ec2d86",
   235 => x"ec2d86ec",
   236 => x"2d86ec2d",
   237 => x"86ec2d86",
   238 => x"ec2d86ec",
   239 => x"2d86ec2d",
   240 => x"86ec2d86",
   241 => x"ec2d86ec",
   242 => x"2d86ec2d",
   243 => x"86ec2d86",
   244 => x"ec2d86ec",
   245 => x"2d86ec2d",
   246 => x"86ec2d86",
   247 => x"ec2d86ec",
   248 => x"2d86ec2d",
   249 => x"86ec2d86",
   250 => x"ec2d86ec",
   251 => x"2d86ec2d",
   252 => x"86ec2d86",
   253 => x"ec2d86ec",
   254 => x"2d86ec2d",
   255 => x"86ec2d86",
   256 => x"ec2d86ec",
   257 => x"2d86ec2d",
   258 => x"86ec2d86",
   259 => x"ec2d86ec",
   260 => x"2d86ec2d",
   261 => x"86ec2d86",
   262 => x"ec2d86ec",
   263 => x"2d86ec2d",
   264 => x"86ec2d86",
   265 => x"ec2d86ec",
   266 => x"2d86ec2d",
   267 => x"86ec2d86",
   268 => x"ec2d86ec",
   269 => x"2d86ec2d",
   270 => x"86ec2d86",
   271 => x"ec2d86ec",
   272 => x"2d86ec2d",
   273 => x"86ec2d86",
   274 => x"ec2d86ec",
   275 => x"2d86ec2d",
   276 => x"86ec2d86",
   277 => x"ec2d86ec",
   278 => x"2d86ec2d",
   279 => x"86ec2d86",
   280 => x"ec2d86ec",
   281 => x"2d86ec2d",
   282 => x"86ec2d86",
   283 => x"ec2d86ec",
   284 => x"2d86ec2d",
   285 => x"86ec2d86",
   286 => x"ec2d86ec",
   287 => x"2d86ec2d",
   288 => x"86ec2d86",
   289 => x"ec2d86ec",
   290 => x"2d86ec2d",
   291 => x"86ec2d86",
   292 => x"ec2d86ec",
   293 => x"2d86ec2d",
   294 => x"86ec2d86",
   295 => x"ec2d86ec",
   296 => x"2d86ec2d",
   297 => x"86ec2d86",
   298 => x"ec2d86ec",
   299 => x"2d86ec2d",
   300 => x"86ec2d86",
   301 => x"ec2d86ec",
   302 => x"2d86ec2d",
   303 => x"86ec2d86",
   304 => x"ec2d86ec",
   305 => x"2d86ec2d",
   306 => x"86ec2d86",
   307 => x"ec2d86ec",
   308 => x"2d86ec2d",
   309 => x"86ec2d86",
   310 => x"ec2d86ec",
   311 => x"2d86ec2d",
   312 => x"86ec2d86",
   313 => x"ec2d86ec",
   314 => x"2d86ec2d",
   315 => x"86ec2d86",
   316 => x"ec2d86ec",
   317 => x"2d86ec2d",
   318 => x"86ec2d86",
   319 => x"ec2d86ec",
   320 => x"2d86ec2d",
   321 => x"86ec2d86",
   322 => x"ec2d86ec",
   323 => x"2d86ec2d",
   324 => x"86ec2d86",
   325 => x"ec2d86ec",
   326 => x"2d86ec2d",
   327 => x"86ec2d86",
   328 => x"ec2d86ec",
   329 => x"2d86ec2d",
   330 => x"86ec2d86",
   331 => x"ec2d86ec",
   332 => x"2d86ec2d",
   333 => x"86ec2d86",
   334 => x"ec2d86ec",
   335 => x"2d86ec2d",
   336 => x"86ec2d86",
   337 => x"ec2d86ec",
   338 => x"2d86ec2d",
   339 => x"86ec2d86",
   340 => x"ec2d86ec",
   341 => x"2d86ec2d",
   342 => x"86ec2d86",
   343 => x"ec2d86ec",
   344 => x"2d86ec2d",
   345 => x"86ec2d86",
   346 => x"ec2d86ec",
   347 => x"2d86ec2d",
   348 => x"86ec2d86",
   349 => x"ec2d86ec",
   350 => x"2d86ec2d",
   351 => x"86ec2d86",
   352 => x"ec2d86ec",
   353 => x"2d86ec2d",
   354 => x"86ec2d86",
   355 => x"ec2d86ec",
   356 => x"2d86ec2d",
   357 => x"86ec2d86",
   358 => x"ec2d86ec",
   359 => x"2d86ec2d",
   360 => x"86ec2d86",
   361 => x"ec2d86ec",
   362 => x"2d86ec2d",
   363 => x"86ec2d86",
   364 => x"ec2d86ec",
   365 => x"2d86ec2d",
   366 => x"86ec2d86",
   367 => x"ec2d86ec",
   368 => x"2d86ec2d",
   369 => x"86ec2d86",
   370 => x"ec2d86ec",
   371 => x"2d86ec2d",
   372 => x"86ec2d86",
   373 => x"ec2d86ec",
   374 => x"2d86ec2d",
   375 => x"86ec2d86",
   376 => x"ec2d86ec",
   377 => x"2d86ec2d",
   378 => x"86ec2d86",
   379 => x"ec2d86ec",
   380 => x"2d86ec2d",
   381 => x"86ec2d86",
   382 => x"ec2d86ec",
   383 => x"2d86ec2d",
   384 => x"86ec2d86",
   385 => x"ec2d86ec",
   386 => x"2d86ec2d",
   387 => x"86ec2d86",
   388 => x"ec2d86ec",
   389 => x"2d86ec2d",
   390 => x"86ec2d86",
   391 => x"ec2d86ec",
   392 => x"2d86ec2d",
   393 => x"86ec2d86",
   394 => x"ec2d86ec",
   395 => x"2d86ec2d",
   396 => x"86ec2d86",
   397 => x"ec2d86ec",
   398 => x"2d86ec2d",
   399 => x"86ec2d86",
   400 => x"ec2d86ec",
   401 => x"2d86ec2d",
   402 => x"86ec2d86",
   403 => x"ec2d86ec",
   404 => x"2d86ec2d",
   405 => x"86ec2d86",
   406 => x"ec2d86ec",
   407 => x"2d86ec2d",
   408 => x"86ec2d86",
   409 => x"ec2d86ec",
   410 => x"2d86ec2d",
   411 => x"86ec2d86",
   412 => x"ec2d86ec",
   413 => x"2d86ec2d",
   414 => x"86ec2d86",
   415 => x"ec2d86ec",
   416 => x"2d86ec2d",
   417 => x"86ec2d86",
   418 => x"ec2d86ec",
   419 => x"2d86ec2d",
   420 => x"86ec2d86",
   421 => x"ec2d86ec",
   422 => x"2d86ec2d",
   423 => x"86ec2d86",
   424 => x"ec2d86ec",
   425 => x"2d86ec2d",
   426 => x"86ec2d86",
   427 => x"ec2d86ec",
   428 => x"2d86ec2d",
   429 => x"86ec2d86",
   430 => x"ec2d86ec",
   431 => x"2d86ec2d",
   432 => x"86ec2d86",
   433 => x"ec2d86ec",
   434 => x"2d86ec2d",
   435 => x"86ec2d86",
   436 => x"ec2d86ec",
   437 => x"2d86ec2d",
   438 => x"86ec2d86",
   439 => x"ec2d86ec",
   440 => x"2d86ec2d",
   441 => x"86ec2d86",
   442 => x"ec2d86ec",
   443 => x"2d86ec2d",
   444 => x"86ec2d86",
   445 => x"ec2d86ec",
   446 => x"2d86ec2d",
   447 => x"86ec2d86",
   448 => x"ec2d86ec",
   449 => x"2d86ec2d",
   450 => x"86ec2d86",
   451 => x"ec2d86ec",
   452 => x"2d86ec2d",
   453 => x"86ec2d86",
   454 => x"ec2d86ec",
   455 => x"2d86ec2d",
   456 => x"86ec2d86",
   457 => x"ec2d86ec",
   458 => x"2d86ec2d",
   459 => x"86ec2d86",
   460 => x"ec2d86ec",
   461 => x"2d86ec2d",
   462 => x"86ec2d86",
   463 => x"ec2d86ec",
   464 => x"2d86ec2d",
   465 => x"86ec2d86",
   466 => x"ec2d86ec",
   467 => x"2d86ec2d",
   468 => x"86ec2d86",
   469 => x"ec2d86ec",
   470 => x"2d86ec2d",
   471 => x"86ec2d86",
   472 => x"ec2d86ec",
   473 => x"2d86ec2d",
   474 => x"86ec2d86",
   475 => x"ec2d86ec",
   476 => x"2d86ec2d",
   477 => x"86ec2d86",
   478 => x"ec2d86ec",
   479 => x"2d86ec2d",
   480 => x"86ec2d86",
   481 => x"ec2d86ec",
   482 => x"2d86ec2d",
   483 => x"86ec2d86",
   484 => x"ec2d86ec",
   485 => x"2d86ec2d",
   486 => x"86ec2d86",
   487 => x"ec2d86ec",
   488 => x"2d86ec2d",
   489 => x"86ec2d86",
   490 => x"ec2d86ec",
   491 => x"2d86ec2d",
   492 => x"86ec2d86",
   493 => x"ec2d86ec",
   494 => x"2d86ec2d",
   495 => x"86ec2d86",
   496 => x"ec2d86ec",
   497 => x"2d86ec2d",
   498 => x"86ec2d86",
   499 => x"ec2d86ec",
   500 => x"2d86ec2d",
   501 => x"86ec2d86",
   502 => x"ec2d86ec",
   503 => x"2d86ec2d",
   504 => x"86ec2d86",
   505 => x"ec2d86ec",
   506 => x"2d86ec2d",
   507 => x"86ec2d86",
   508 => x"ec2d86ec",
   509 => x"2d86ec2d",
   510 => x"86ec2d86",
   511 => x"ec2d86ec",
   512 => x"2d86ec2d",
   513 => x"86ec2d86",
   514 => x"ec2d86ec",
   515 => x"2d86ec2d",
   516 => x"86ec2d86",
   517 => x"ec2d86ec",
   518 => x"2d86ec2d",
   519 => x"86ec2d86",
   520 => x"ec2d86ec",
   521 => x"2d86ec2d",
   522 => x"86ec2d86",
   523 => x"ec2d86ec",
   524 => x"2d86ec2d",
   525 => x"86ec2d86",
   526 => x"ec2d86ec",
   527 => x"2d86ec2d",
   528 => x"86ec2d86",
   529 => x"ec2d86ec",
   530 => x"2d86ec2d",
   531 => x"86ec2d86",
   532 => x"ec2d86ec",
   533 => x"2d86ec2d",
   534 => x"86ec2d86",
   535 => x"ec2d86ec",
   536 => x"2d86ec2d",
   537 => x"86ec2d86",
   538 => x"ec2d86ec",
   539 => x"2d86ec2d",
   540 => x"86ec2d86",
   541 => x"ec2d86ec",
   542 => x"2d86ec2d",
   543 => x"86ec2d86",
   544 => x"ec2d86ec",
   545 => x"2d86ec2d",
   546 => x"86ec2d86",
   547 => x"ec2d86ec",
   548 => x"2d86ec2d",
   549 => x"86ec2d86",
   550 => x"ec2d86ec",
   551 => x"2d86ec2d",
   552 => x"86ec2d86",
   553 => x"ec2d86ec",
   554 => x"2d86ec2d",
   555 => x"86ec2d86",
   556 => x"ec2d86ec",
   557 => x"2d86ec2d",
   558 => x"86ec2d86",
   559 => x"ec2d86ec",
   560 => x"2d86ec2d",
   561 => x"86ec2d86",
   562 => x"ec2d86ec",
   563 => x"2d86ec2d",
   564 => x"86ec2d86",
   565 => x"ec2d86ec",
   566 => x"2d86ec2d",
   567 => x"86ec2d86",
   568 => x"ec2d86ec",
   569 => x"2d86ec2d",
   570 => x"86ec2d86",
   571 => x"ec2d86ec",
   572 => x"2d86ec2d",
   573 => x"86ec2d86",
   574 => x"ec2d86ec",
   575 => x"2d86ec2d",
   576 => x"86ec2d86",
   577 => x"ec2d86ec",
   578 => x"2d86ec2d",
   579 => x"86ec2d86",
   580 => x"ec2d86ec",
   581 => x"2d86ec2d",
   582 => x"86ec2d86",
   583 => x"ec2d86ec",
   584 => x"2d86ec2d",
   585 => x"86ec2d86",
   586 => x"ec2d86ec",
   587 => x"2d86ec2d",
   588 => x"86ec2d86",
   589 => x"ec2d86ec",
   590 => x"2d86ec2d",
   591 => x"86ec2d86",
   592 => x"ec2d86ec",
   593 => x"2d86ec2d",
   594 => x"86ec2d86",
   595 => x"ec2d86ec",
   596 => x"2d86ec2d",
   597 => x"86ec2d86",
   598 => x"ec2d86ec",
   599 => x"2d86ec2d",
   600 => x"86ec2d86",
   601 => x"ec2d86ec",
   602 => x"2d86ec2d",
   603 => x"86ec2d86",
   604 => x"ec2d86ec",
   605 => x"2d86ec2d",
   606 => x"86ec2d86",
   607 => x"ec2d86ec",
   608 => x"2d86ec2d",
   609 => x"86ec2d86",
   610 => x"ec2d86ec",
   611 => x"2d86ec2d",
   612 => x"86ec2d86",
   613 => x"ec2d86ec",
   614 => x"2d86ec2d",
   615 => x"86ec2d86",
   616 => x"ec2d86ec",
   617 => x"2d86ec2d",
   618 => x"86ec2d86",
   619 => x"ec2d86ec",
   620 => x"2d86ec2d",
   621 => x"86ec2d86",
   622 => x"ec2d86ec",
   623 => x"2d86ec2d",
   624 => x"86ec2d86",
   625 => x"ec2d86ec",
   626 => x"2d86ec2d",
   627 => x"86ec2d86",
   628 => x"ec2d86ec",
   629 => x"2d86ec2d",
   630 => x"86ec2d86",
   631 => x"ec2d86ec",
   632 => x"2d86ec2d",
   633 => x"86ec2d86",
   634 => x"ec2d86ec",
   635 => x"2d86ec2d",
   636 => x"86ec2d86",
   637 => x"ec2d86ec",
   638 => x"2d86ec2d",
   639 => x"86ec2d86",
   640 => x"ec2d86ec",
   641 => x"2d86ec2d",
   642 => x"86ec2d86",
   643 => x"ec2d86ec",
   644 => x"2d86ec2d",
   645 => x"86ec2d86",
   646 => x"ec2d86ec",
   647 => x"2d86ec2d",
   648 => x"86ec2d86",
   649 => x"ec2d86ec",
   650 => x"2d86ec2d",
   651 => x"86ec2d86",
   652 => x"ec2d86ec",
   653 => x"2d86ec2d",
   654 => x"86ec2d86",
   655 => x"ec2d86ec",
   656 => x"2d86ec2d",
   657 => x"86ec2d86",
   658 => x"ec2d86ec",
   659 => x"2d86ec2d",
   660 => x"86ec2d04",
   661 => x"0402dc05",
   662 => x"0d7a5380",
   663 => x"59840bec",
   664 => x"0c725280",
   665 => x"d3b451bf",
   666 => x"ee2d80d3",
   667 => x"9808792e",
   668 => x"81c43880",
   669 => x"d3b80855",
   670 => x"74852e09",
   671 => x"8106bb38",
   672 => x"725186c5",
   673 => x"2d87932d",
   674 => x"87932d87",
   675 => x"932d8793",
   676 => x"2d87932d",
   677 => x"87932d80",
   678 => x"d3e80888",
   679 => x"2a708106",
   680 => x"51537279",
   681 => x"2e883880",
   682 => x"cfb05195",
   683 => x"b20480ce",
   684 => x"a051a191",
   685 => x"2d815396",
   686 => x"e70474f8",
   687 => x"0ca50bec",
   688 => x"0c87932d",
   689 => x"840bec0c",
   690 => x"78ff1655",
   691 => x"5873802e",
   692 => x"8b388118",
   693 => x"74812a55",
   694 => x"5895cd04",
   695 => x"f7185881",
   696 => x"59807525",
   697 => x"80d03877",
   698 => x"52735184",
   699 => x"a82d80d4",
   700 => x"885280d3",
   701 => x"b45180c2",
   702 => x"c02d80d3",
   703 => x"9808802e",
   704 => x"9b3880d4",
   705 => x"885783fc",
   706 => x"56767084",
   707 => x"055808e8",
   708 => x"0cfc1656",
   709 => x"758025f1",
   710 => x"3896a404",
   711 => x"80d39808",
   712 => x"59848055",
   713 => x"80d3b451",
   714 => x"80c2902d",
   715 => x"fc801581",
   716 => x"15555595",
   717 => x"e1048051",
   718 => x"86ff2d78",
   719 => x"802e9f38",
   720 => x"80d3e808",
   721 => x"882a7081",
   722 => x"06515372",
   723 => x"802e8838",
   724 => x"80cfb051",
   725 => x"96e20480",
   726 => x"cea05196",
   727 => x"e20480d0",
   728 => x"c051a191",
   729 => x"2d785372",
   730 => x"80d3980c",
   731 => x"02a4050d",
   732 => x"0402e805",
   733 => x"0d805186",
   734 => x"ff2d840b",
   735 => x"ec0c9ea9",
   736 => x"2d9ad42d",
   737 => x"81f92d83",
   738 => x"539e8c2d",
   739 => x"8151858d",
   740 => x"2dff1353",
   741 => x"728025f1",
   742 => x"38840bec",
   743 => x"0c80ccd0",
   744 => x"5186c52d",
   745 => x"b6a32d80",
   746 => x"d3980880",
   747 => x"2e838e38",
   748 => x"810bec0c",
   749 => x"840bec0c",
   750 => x"80c9a852",
   751 => x"80d3b451",
   752 => x"bfee2d80",
   753 => x"d3980880",
   754 => x"2e80cc38",
   755 => x"80d48852",
   756 => x"80d3b451",
   757 => x"80c2c02d",
   758 => x"80d39808",
   759 => x"802eb838",
   760 => x"80d4880b",
   761 => x"80f52d80",
   762 => x"d1c40c80",
   763 => x"d4890b80",
   764 => x"f52d80d1",
   765 => x"c80c80d4",
   766 => x"8a0b80f5",
   767 => x"2d80d1cc",
   768 => x"0c80d48b",
   769 => x"0b80f52d",
   770 => x"80d1d00c",
   771 => x"80d48c0b",
   772 => x"80f52d80",
   773 => x"d1d40c80",
   774 => x"c9b85280",
   775 => x"d3b451bf",
   776 => x"ee2d80d3",
   777 => x"9808802e",
   778 => x"80cc3880",
   779 => x"d4885280",
   780 => x"d3b45180",
   781 => x"c2c02d80",
   782 => x"d3980880",
   783 => x"2eb83880",
   784 => x"d4880b80",
   785 => x"f52d80d1",
   786 => x"b00c80d4",
   787 => x"890b80f5",
   788 => x"2d80d1b4",
   789 => x"0c80d48a",
   790 => x"0b80f52d",
   791 => x"80d1b80c",
   792 => x"80d48b0b",
   793 => x"80f52d80",
   794 => x"d1bc0c80",
   795 => x"d48c0b80",
   796 => x"f52d80d1",
   797 => x"c00c94d5",
   798 => x"5180c992",
   799 => x"2d900b80",
   800 => x"d1ac0c90",
   801 => x"0bfc0c80",
   802 => x"d3e80888",
   803 => x"2a708106",
   804 => x"51537280",
   805 => x"2e883880",
   806 => x"cfb05199",
   807 => x"a20480ce",
   808 => x"a051a191",
   809 => x"2d850b80",
   810 => x"d3fc0c9e",
   811 => x"e22d9ae0",
   812 => x"2da1a42d",
   813 => x"80d39808",
   814 => x"80d3e808",
   815 => x"882a7081",
   816 => x"06515456",
   817 => x"72802eaa",
   818 => x"3880d080",
   819 => x"0b80f52d",
   820 => x"80d08c0b",
   821 => x"80f52d71",
   822 => x"842b7185",
   823 => x"2b0780d0",
   824 => x"980b80f5",
   825 => x"2d70822b",
   826 => x"72075253",
   827 => x"5656539a",
   828 => x"8a0480ce",
   829 => x"f00b80f5",
   830 => x"2d80cefc",
   831 => x"0b80f52d",
   832 => x"71842b71",
   833 => x"852b0756",
   834 => x"545580d1",
   835 => x"ac087081",
   836 => x"06545572",
   837 => x"802e8538",
   838 => x"73810754",
   839 => x"74812a70",
   840 => x"81065153",
   841 => x"72802e85",
   842 => x"38738207",
   843 => x"5473fc0c",
   844 => x"86537583",
   845 => x"38845372",
   846 => x"ec0c99ae",
   847 => x"04800b80",
   848 => x"d3980c02",
   849 => x"98050d04",
   850 => x"71980c04",
   851 => x"ffb00880",
   852 => x"d3980c04",
   853 => x"810bffb0",
   854 => x"0c04800b",
   855 => x"ffb00c04",
   856 => x"02f4050d",
   857 => x"9bee0480",
   858 => x"d3980881",
   859 => x"f02e0981",
   860 => x"068a3881",
   861 => x"0b80d1a4",
   862 => x"0c9bee04",
   863 => x"80d39808",
   864 => x"81e02e09",
   865 => x"81068a38",
   866 => x"810b80d1",
   867 => x"a80c9bee",
   868 => x"0480d398",
   869 => x"085280d1",
   870 => x"a808802e",
   871 => x"893880d3",
   872 => x"98088180",
   873 => x"05527184",
   874 => x"2c728f06",
   875 => x"535380d1",
   876 => x"a408802e",
   877 => x"9a387284",
   878 => x"2980d0e4",
   879 => x"05721381",
   880 => x"712b7009",
   881 => x"73080673",
   882 => x"0c515353",
   883 => x"9be20472",
   884 => x"842980d0",
   885 => x"e4057213",
   886 => x"83712b72",
   887 => x"0807720c",
   888 => x"5353800b",
   889 => x"80d1a80c",
   890 => x"800b80d1",
   891 => x"a40c80d3",
   892 => x"c0519cf5",
   893 => x"2d80d398",
   894 => x"08ff24fe",
   895 => x"ea38800b",
   896 => x"80d3980c",
   897 => x"028c050d",
   898 => x"0402f805",
   899 => x"0d80d0e4",
   900 => x"528f5180",
   901 => x"72708405",
   902 => x"540cff11",
   903 => x"51708025",
   904 => x"f2380288",
   905 => x"050d0402",
   906 => x"f0050d75",
   907 => x"519ada2d",
   908 => x"70822cfc",
   909 => x"0680d0e4",
   910 => x"1172109e",
   911 => x"06710870",
   912 => x"722a7083",
   913 => x"0682742b",
   914 => x"70097406",
   915 => x"760c5451",
   916 => x"56575351",
   917 => x"539ad42d",
   918 => x"7180d398",
   919 => x"0c029005",
   920 => x"0d0402fc",
   921 => x"050d7251",
   922 => x"80710c80",
   923 => x"0b84120c",
   924 => x"0284050d",
   925 => x"0402f005",
   926 => x"0d757008",
   927 => x"84120853",
   928 => x"5353ff54",
   929 => x"71712ea8",
   930 => x"389ada2d",
   931 => x"84130870",
   932 => x"84291488",
   933 => x"11700870",
   934 => x"81ff0684",
   935 => x"18088111",
   936 => x"8706841a",
   937 => x"0c535155",
   938 => x"5151519a",
   939 => x"d42d7154",
   940 => x"7380d398",
   941 => x"0c029005",
   942 => x"0d0402f4",
   943 => x"050d9ada",
   944 => x"2de00870",
   945 => x"8b2a7081",
   946 => x"06515253",
   947 => x"70802ea1",
   948 => x"3880d3c0",
   949 => x"08708429",
   950 => x"80d3c805",
   951 => x"7481ff06",
   952 => x"710c5151",
   953 => x"80d3c008",
   954 => x"81118706",
   955 => x"80d3c00c",
   956 => x"51728c2c",
   957 => x"83ff0680",
   958 => x"d3e80c80",
   959 => x"0b80d3ec",
   960 => x"0c9acc2d",
   961 => x"9ad42d02",
   962 => x"8c050d04",
   963 => x"02fc050d",
   964 => x"9ada2d81",
   965 => x"0b80d3ec",
   966 => x"0c9ad42d",
   967 => x"80d3ec08",
   968 => x"5170f938",
   969 => x"0284050d",
   970 => x"0402fc05",
   971 => x"0d80d3c0",
   972 => x"519ce22d",
   973 => x"9c892d9d",
   974 => x"ba519ac8",
   975 => x"2d028405",
   976 => x"0d0402fc",
   977 => x"050d8fcf",
   978 => x"5186ec2d",
   979 => x"ff115170",
   980 => x"8025f638",
   981 => x"0284050d",
   982 => x"0480d3f4",
   983 => x"0880d398",
   984 => x"0c0402fc",
   985 => x"050d810b",
   986 => x"80d1d80c",
   987 => x"8151858d",
   988 => x"2d028405",
   989 => x"0d0402fc",
   990 => x"050d9f80",
   991 => x"049ae02d",
   992 => x"80f6519c",
   993 => x"a72d80d3",
   994 => x"9808f238",
   995 => x"80da519c",
   996 => x"a72d80d3",
   997 => x"9808e638",
   998 => x"80d1d408",
   999 => x"519ca72d",
  1000 => x"80d39808",
  1001 => x"d83880d3",
  1002 => x"980880d1",
  1003 => x"d80c80d3",
  1004 => x"98085185",
  1005 => x"8d2d0284",
  1006 => x"050d0402",
  1007 => x"ec050d76",
  1008 => x"54805287",
  1009 => x"0b881580",
  1010 => x"f52d5653",
  1011 => x"74722483",
  1012 => x"38a05372",
  1013 => x"5183842d",
  1014 => x"81128b15",
  1015 => x"80f52d54",
  1016 => x"52727225",
  1017 => x"de380294",
  1018 => x"050d0402",
  1019 => x"f0050d80",
  1020 => x"d3f40854",
  1021 => x"81f92d80",
  1022 => x"0b80d3f8",
  1023 => x"0c730880",
  1024 => x"2e818938",
  1025 => x"820b80d3",
  1026 => x"ac0c80d3",
  1027 => x"f8088f06",
  1028 => x"80d3a80c",
  1029 => x"73085271",
  1030 => x"832e9638",
  1031 => x"71832689",
  1032 => x"3871812e",
  1033 => x"b038a0f5",
  1034 => x"0471852e",
  1035 => x"a038a0f5",
  1036 => x"04881480",
  1037 => x"f52d8415",
  1038 => x"0880cce8",
  1039 => x"53545286",
  1040 => x"c52d7184",
  1041 => x"29137008",
  1042 => x"5252a0f9",
  1043 => x"0473519f",
  1044 => x"bb2da0f5",
  1045 => x"0480d1ac",
  1046 => x"08881508",
  1047 => x"2c708106",
  1048 => x"51527180",
  1049 => x"2e883880",
  1050 => x"ccec51a0",
  1051 => x"f20480cc",
  1052 => x"f05186c5",
  1053 => x"2d841408",
  1054 => x"5186c52d",
  1055 => x"80d3f808",
  1056 => x"810580d3",
  1057 => x"f80c8c14",
  1058 => x"549ffd04",
  1059 => x"0290050d",
  1060 => x"047180d3",
  1061 => x"f40c9feb",
  1062 => x"2d80d3f8",
  1063 => x"08ff0580",
  1064 => x"d3fc0c04",
  1065 => x"02e8050d",
  1066 => x"80d3f408",
  1067 => x"80d48008",
  1068 => x"575580f6",
  1069 => x"519ca72d",
  1070 => x"80d39808",
  1071 => x"812a7081",
  1072 => x"06515271",
  1073 => x"802ea238",
  1074 => x"a1ce049a",
  1075 => x"e02d80f6",
  1076 => x"519ca72d",
  1077 => x"80d39808",
  1078 => x"f23880d1",
  1079 => x"d8088132",
  1080 => x"7080d1d8",
  1081 => x"0c51858d",
  1082 => x"2d800b80",
  1083 => x"d3f00c8c",
  1084 => x"519ca72d",
  1085 => x"80d39808",
  1086 => x"812a7081",
  1087 => x"06515271",
  1088 => x"802e80d1",
  1089 => x"3880d1b0",
  1090 => x"0880d1c4",
  1091 => x"0880d1b0",
  1092 => x"0c80d1c4",
  1093 => x"0c80d1b4",
  1094 => x"0880d1c8",
  1095 => x"0880d1b4",
  1096 => x"0c80d1c8",
  1097 => x"0c80d1b8",
  1098 => x"0880d1cc",
  1099 => x"0880d1b8",
  1100 => x"0c80d1cc",
  1101 => x"0c80d1bc",
  1102 => x"0880d1d0",
  1103 => x"0880d1bc",
  1104 => x"0c80d1d0",
  1105 => x"0c80d1c0",
  1106 => x"0880d1d4",
  1107 => x"0880d1c0",
  1108 => x"0c80d1d4",
  1109 => x"0c80d3e8",
  1110 => x"08a00652",
  1111 => x"80722596",
  1112 => x"389ec22d",
  1113 => x"9ae02d80",
  1114 => x"d1d80881",
  1115 => x"327080d1",
  1116 => x"d80c5185",
  1117 => x"8d2d80d1",
  1118 => x"d80882ef",
  1119 => x"3880d1c4",
  1120 => x"08519ca7",
  1121 => x"2d80d398",
  1122 => x"08802e8b",
  1123 => x"3880d3f0",
  1124 => x"08810780",
  1125 => x"d3f00c80",
  1126 => x"d1c80851",
  1127 => x"9ca72d80",
  1128 => x"d3980880",
  1129 => x"2e8b3880",
  1130 => x"d3f00882",
  1131 => x"0780d3f0",
  1132 => x"0c80d1cc",
  1133 => x"08519ca7",
  1134 => x"2d80d398",
  1135 => x"08802e8b",
  1136 => x"3880d3f0",
  1137 => x"08840780",
  1138 => x"d3f00c80",
  1139 => x"d1d00851",
  1140 => x"9ca72d80",
  1141 => x"d3980880",
  1142 => x"2e8b3880",
  1143 => x"d3f00888",
  1144 => x"0780d3f0",
  1145 => x"0c80d1d4",
  1146 => x"08519ca7",
  1147 => x"2d80d398",
  1148 => x"08802e8b",
  1149 => x"3880d3f0",
  1150 => x"08900780",
  1151 => x"d3f00c80",
  1152 => x"d1b00851",
  1153 => x"9ca72d80",
  1154 => x"d3980880",
  1155 => x"2e8c3880",
  1156 => x"d3f00882",
  1157 => x"800780d3",
  1158 => x"f00c80d1",
  1159 => x"b408519c",
  1160 => x"a72d80d3",
  1161 => x"9808802e",
  1162 => x"8c3880d3",
  1163 => x"f0088480",
  1164 => x"0780d3f0",
  1165 => x"0c80d1b8",
  1166 => x"08519ca7",
  1167 => x"2d80d398",
  1168 => x"08802e8c",
  1169 => x"3880d3f0",
  1170 => x"08888007",
  1171 => x"80d3f00c",
  1172 => x"80d1bc08",
  1173 => x"519ca72d",
  1174 => x"80d39808",
  1175 => x"802e8c38",
  1176 => x"80d3f008",
  1177 => x"90800780",
  1178 => x"d3f00c80",
  1179 => x"d1c00851",
  1180 => x"9ca72d80",
  1181 => x"d3980880",
  1182 => x"2e8c3880",
  1183 => x"d3f008a0",
  1184 => x"800780d3",
  1185 => x"f00c9451",
  1186 => x"9ca72d80",
  1187 => x"d3980852",
  1188 => x"91519ca7",
  1189 => x"2d7180d3",
  1190 => x"98080652",
  1191 => x"80e6519c",
  1192 => x"a72d7180",
  1193 => x"d3980806",
  1194 => x"5271802e",
  1195 => x"8d3880d3",
  1196 => x"f0088480",
  1197 => x"800780d3",
  1198 => x"f00c80fe",
  1199 => x"519ca72d",
  1200 => x"80d39808",
  1201 => x"5287519c",
  1202 => x"a72d7180",
  1203 => x"d3980807",
  1204 => x"5271802e",
  1205 => x"8d3880d3",
  1206 => x"f0088880",
  1207 => x"800780d3",
  1208 => x"f00c80d3",
  1209 => x"f008ed0c",
  1210 => x"adf60494",
  1211 => x"519ca72d",
  1212 => x"80d39808",
  1213 => x"5291519c",
  1214 => x"a72d7180",
  1215 => x"d3980806",
  1216 => x"5280e651",
  1217 => x"9ca72d71",
  1218 => x"80d39808",
  1219 => x"06527180",
  1220 => x"2e8d3880",
  1221 => x"d3f00884",
  1222 => x"80800780",
  1223 => x"d3f00c80",
  1224 => x"fe519ca7",
  1225 => x"2d80d398",
  1226 => x"08528751",
  1227 => x"9ca72d71",
  1228 => x"80d39808",
  1229 => x"07527180",
  1230 => x"2e8d3880",
  1231 => x"d3f00888",
  1232 => x"80800780",
  1233 => x"d3f00c80",
  1234 => x"d3f008ed",
  1235 => x"0c81f551",
  1236 => x"9ca72d80",
  1237 => x"d3980881",
  1238 => x"2a708106",
  1239 => x"515271a4",
  1240 => x"3880d1c4",
  1241 => x"08519ca7",
  1242 => x"2d80d398",
  1243 => x"08812a70",
  1244 => x"81065152",
  1245 => x"718e3880",
  1246 => x"d3e80881",
  1247 => x"06528072",
  1248 => x"2580c238",
  1249 => x"80d3e808",
  1250 => x"81065280",
  1251 => x"72258438",
  1252 => x"9ec22d80",
  1253 => x"d3fc0852",
  1254 => x"71802e8a",
  1255 => x"38ff1280",
  1256 => x"d3fc0ca7",
  1257 => x"c50480d3",
  1258 => x"f8081080",
  1259 => x"d3f80805",
  1260 => x"70842916",
  1261 => x"51528812",
  1262 => x"08802e89",
  1263 => x"38ff5188",
  1264 => x"12085271",
  1265 => x"2d81f251",
  1266 => x"9ca72d80",
  1267 => x"d3980881",
  1268 => x"2a708106",
  1269 => x"515271a4",
  1270 => x"3880d1c8",
  1271 => x"08519ca7",
  1272 => x"2d80d398",
  1273 => x"08812a70",
  1274 => x"81065152",
  1275 => x"718e3880",
  1276 => x"d3e80882",
  1277 => x"06528072",
  1278 => x"2580c338",
  1279 => x"80d3e808",
  1280 => x"82065280",
  1281 => x"72258438",
  1282 => x"9ec22d80",
  1283 => x"d3f808ff",
  1284 => x"1180d3fc",
  1285 => x"08565353",
  1286 => x"7372258a",
  1287 => x"38811480",
  1288 => x"d3fc0ca8",
  1289 => x"be047210",
  1290 => x"13708429",
  1291 => x"16515288",
  1292 => x"1208802e",
  1293 => x"8938fe51",
  1294 => x"88120852",
  1295 => x"712d81fd",
  1296 => x"519ca72d",
  1297 => x"80d39808",
  1298 => x"812a7081",
  1299 => x"06515271",
  1300 => x"a43880d1",
  1301 => x"cc08519c",
  1302 => x"a72d80d3",
  1303 => x"9808812a",
  1304 => x"70810651",
  1305 => x"52718e38",
  1306 => x"80d3e808",
  1307 => x"84065280",
  1308 => x"722580c0",
  1309 => x"3880d3e8",
  1310 => x"08840652",
  1311 => x"80722584",
  1312 => x"389ec22d",
  1313 => x"80d3fc08",
  1314 => x"802e8a38",
  1315 => x"800b80d3",
  1316 => x"fc0ca9b4",
  1317 => x"0480d3f8",
  1318 => x"081080d3",
  1319 => x"f8080570",
  1320 => x"84291651",
  1321 => x"52881208",
  1322 => x"802e8938",
  1323 => x"fd518812",
  1324 => x"0852712d",
  1325 => x"81fa519c",
  1326 => x"a72d80d3",
  1327 => x"9808812a",
  1328 => x"70810651",
  1329 => x"5271a438",
  1330 => x"80d1d008",
  1331 => x"519ca72d",
  1332 => x"80d39808",
  1333 => x"812a7081",
  1334 => x"06515271",
  1335 => x"8e3880d3",
  1336 => x"e8088806",
  1337 => x"52807225",
  1338 => x"80c03880",
  1339 => x"d3e80888",
  1340 => x"06528072",
  1341 => x"2584389e",
  1342 => x"c22d80d3",
  1343 => x"f808ff11",
  1344 => x"545280d3",
  1345 => x"fc087325",
  1346 => x"89387280",
  1347 => x"d3fc0caa",
  1348 => x"aa047110",
  1349 => x"12708429",
  1350 => x"16515288",
  1351 => x"1208802e",
  1352 => x"8938fc51",
  1353 => x"88120852",
  1354 => x"712d80d3",
  1355 => x"fc087053",
  1356 => x"5473802e",
  1357 => x"8a388c15",
  1358 => x"ff155555",
  1359 => x"aab10482",
  1360 => x"0b80d3ac",
  1361 => x"0c718f06",
  1362 => x"80d3a80c",
  1363 => x"81eb519c",
  1364 => x"a72d80d3",
  1365 => x"9808812a",
  1366 => x"70810651",
  1367 => x"5271802e",
  1368 => x"ad387408",
  1369 => x"852e0981",
  1370 => x"06a43888",
  1371 => x"1580f52d",
  1372 => x"ff055271",
  1373 => x"881681b7",
  1374 => x"2d71982b",
  1375 => x"52718025",
  1376 => x"8838800b",
  1377 => x"881681b7",
  1378 => x"2d74519f",
  1379 => x"bb2d81f4",
  1380 => x"519ca72d",
  1381 => x"80d39808",
  1382 => x"812a7081",
  1383 => x"06515271",
  1384 => x"802eb338",
  1385 => x"7408852e",
  1386 => x"098106aa",
  1387 => x"38881580",
  1388 => x"f52d8105",
  1389 => x"52718816",
  1390 => x"81b72d71",
  1391 => x"81ff068b",
  1392 => x"1680f52d",
  1393 => x"54527272",
  1394 => x"27873872",
  1395 => x"881681b7",
  1396 => x"2d74519f",
  1397 => x"bb2d80da",
  1398 => x"519ca72d",
  1399 => x"80d39808",
  1400 => x"812a7081",
  1401 => x"06515271",
  1402 => x"8e3880d3",
  1403 => x"e8089006",
  1404 => x"52807225",
  1405 => x"81bc3880",
  1406 => x"d3f40880",
  1407 => x"d3e80890",
  1408 => x"06535380",
  1409 => x"72258438",
  1410 => x"9ec22d80",
  1411 => x"d3fc0854",
  1412 => x"73802e8a",
  1413 => x"388c13ff",
  1414 => x"155553ac",
  1415 => x"90047208",
  1416 => x"5271822e",
  1417 => x"a6387182",
  1418 => x"26893871",
  1419 => x"812eaa38",
  1420 => x"adb20471",
  1421 => x"832eb438",
  1422 => x"71842e09",
  1423 => x"810680f2",
  1424 => x"38881308",
  1425 => x"51a1912d",
  1426 => x"adb20480",
  1427 => x"d3fc0851",
  1428 => x"88130852",
  1429 => x"712dadb2",
  1430 => x"04810b88",
  1431 => x"14082b80",
  1432 => x"d1ac0832",
  1433 => x"80d1ac0c",
  1434 => x"ad860488",
  1435 => x"1380f52d",
  1436 => x"81058b14",
  1437 => x"80f52d53",
  1438 => x"54717424",
  1439 => x"83388054",
  1440 => x"73881481",
  1441 => x"b72d9feb",
  1442 => x"2dadb204",
  1443 => x"7508802e",
  1444 => x"a4387508",
  1445 => x"519ca72d",
  1446 => x"80d39808",
  1447 => x"81065271",
  1448 => x"802e8c38",
  1449 => x"80d3fc08",
  1450 => x"51841608",
  1451 => x"52712d88",
  1452 => x"165675d8",
  1453 => x"38805480",
  1454 => x"0b80d3ac",
  1455 => x"0c738f06",
  1456 => x"80d3a80c",
  1457 => x"a0527380",
  1458 => x"d3fc082e",
  1459 => x"09810699",
  1460 => x"3880d3f8",
  1461 => x"08ff0574",
  1462 => x"32700981",
  1463 => x"05707207",
  1464 => x"9f2a9171",
  1465 => x"31515153",
  1466 => x"53715183",
  1467 => x"842d8114",
  1468 => x"548e7425",
  1469 => x"c23880d1",
  1470 => x"d80880d3",
  1471 => x"980c0298",
  1472 => x"050d0402",
  1473 => x"f4050dd4",
  1474 => x"5281ff72",
  1475 => x"0c710853",
  1476 => x"81ff720c",
  1477 => x"72882b83",
  1478 => x"fe800672",
  1479 => x"087081ff",
  1480 => x"06515253",
  1481 => x"81ff720c",
  1482 => x"72710788",
  1483 => x"2b720870",
  1484 => x"81ff0651",
  1485 => x"525381ff",
  1486 => x"720c7271",
  1487 => x"07882b72",
  1488 => x"087081ff",
  1489 => x"06720780",
  1490 => x"d3980c52",
  1491 => x"53028c05",
  1492 => x"0d0402f4",
  1493 => x"050d7476",
  1494 => x"7181ff06",
  1495 => x"d40c5353",
  1496 => x"80d48408",
  1497 => x"85387189",
  1498 => x"2b527198",
  1499 => x"2ad40c71",
  1500 => x"902a7081",
  1501 => x"ff06d40c",
  1502 => x"5171882a",
  1503 => x"7081ff06",
  1504 => x"d40c5171",
  1505 => x"81ff06d4",
  1506 => x"0c72902a",
  1507 => x"7081ff06",
  1508 => x"d40c51d4",
  1509 => x"087081ff",
  1510 => x"06515182",
  1511 => x"b8bf5270",
  1512 => x"81ff2e09",
  1513 => x"81069438",
  1514 => x"81ff0bd4",
  1515 => x"0cd40870",
  1516 => x"81ff06ff",
  1517 => x"14545151",
  1518 => x"71e53870",
  1519 => x"80d3980c",
  1520 => x"028c050d",
  1521 => x"0402fc05",
  1522 => x"0d81c751",
  1523 => x"81ff0bd4",
  1524 => x"0cff1151",
  1525 => x"708025f4",
  1526 => x"38028405",
  1527 => x"0d0402f4",
  1528 => x"050d81ff",
  1529 => x"0bd40c93",
  1530 => x"53805287",
  1531 => x"fc80c151",
  1532 => x"aed22d80",
  1533 => x"d398088b",
  1534 => x"3881ff0b",
  1535 => x"d40c8153",
  1536 => x"b08c04af",
  1537 => x"c52dff13",
  1538 => x"5372de38",
  1539 => x"7280d398",
  1540 => x"0c028c05",
  1541 => x"0d0402ec",
  1542 => x"050d810b",
  1543 => x"80d4840c",
  1544 => x"8454d008",
  1545 => x"708f2a70",
  1546 => x"81065151",
  1547 => x"5372f338",
  1548 => x"72d00caf",
  1549 => x"c52d80cc",
  1550 => x"f45186c5",
  1551 => x"2dd00870",
  1552 => x"8f2a7081",
  1553 => x"06515153",
  1554 => x"72f33881",
  1555 => x"0bd00cb1",
  1556 => x"53805284",
  1557 => x"d480c051",
  1558 => x"aed22d80",
  1559 => x"d3980881",
  1560 => x"2e933872",
  1561 => x"822ebf38",
  1562 => x"ff135372",
  1563 => x"e438ff14",
  1564 => x"5473ffae",
  1565 => x"38afc52d",
  1566 => x"83aa5284",
  1567 => x"9c80c851",
  1568 => x"aed22d80",
  1569 => x"d3980881",
  1570 => x"2e098106",
  1571 => x"9338ae83",
  1572 => x"2d80d398",
  1573 => x"0883ffff",
  1574 => x"06537283",
  1575 => x"aa2e9f38",
  1576 => x"afde2db1",
  1577 => x"b90480cd",
  1578 => x"805186c5",
  1579 => x"2d8053b3",
  1580 => x"8e0480cd",
  1581 => x"985186c5",
  1582 => x"2d8054b2",
  1583 => x"df0481ff",
  1584 => x"0bd40cb1",
  1585 => x"54afc52d",
  1586 => x"8fcf5380",
  1587 => x"5287fc80",
  1588 => x"f751aed2",
  1589 => x"2d80d398",
  1590 => x"085580d3",
  1591 => x"9808812e",
  1592 => x"0981069c",
  1593 => x"3881ff0b",
  1594 => x"d40c820a",
  1595 => x"52849c80",
  1596 => x"e951aed2",
  1597 => x"2d80d398",
  1598 => x"08802e8d",
  1599 => x"38afc52d",
  1600 => x"ff135372",
  1601 => x"c638b2d2",
  1602 => x"0481ff0b",
  1603 => x"d40c80d3",
  1604 => x"98085287",
  1605 => x"fc80fa51",
  1606 => x"aed22d80",
  1607 => x"d39808b2",
  1608 => x"3881ff0b",
  1609 => x"d40cd408",
  1610 => x"5381ff0b",
  1611 => x"d40c81ff",
  1612 => x"0bd40c81",
  1613 => x"ff0bd40c",
  1614 => x"81ff0bd4",
  1615 => x"0c72862a",
  1616 => x"70810676",
  1617 => x"56515372",
  1618 => x"963880d3",
  1619 => x"980854b2",
  1620 => x"df047382",
  1621 => x"2efedb38",
  1622 => x"ff145473",
  1623 => x"fee73873",
  1624 => x"80d4840c",
  1625 => x"738b3881",
  1626 => x"5287fc80",
  1627 => x"d051aed2",
  1628 => x"2d81ff0b",
  1629 => x"d40cd008",
  1630 => x"708f2a70",
  1631 => x"81065151",
  1632 => x"5372f338",
  1633 => x"72d00c81",
  1634 => x"ff0bd40c",
  1635 => x"81537280",
  1636 => x"d3980c02",
  1637 => x"94050d04",
  1638 => x"02e8050d",
  1639 => x"78558056",
  1640 => x"81ff0bd4",
  1641 => x"0cd00870",
  1642 => x"8f2a7081",
  1643 => x"06515153",
  1644 => x"72f33882",
  1645 => x"810bd00c",
  1646 => x"81ff0bd4",
  1647 => x"0c775287",
  1648 => x"fc80d151",
  1649 => x"aed22d80",
  1650 => x"dbc6df54",
  1651 => x"80d39808",
  1652 => x"802e8b38",
  1653 => x"80cdb851",
  1654 => x"86c52db4",
  1655 => x"b20481ff",
  1656 => x"0bd40cd4",
  1657 => x"087081ff",
  1658 => x"06515372",
  1659 => x"81fe2e09",
  1660 => x"81069e38",
  1661 => x"80ff53ae",
  1662 => x"832d80d3",
  1663 => x"98087570",
  1664 => x"8405570c",
  1665 => x"ff135372",
  1666 => x"8025ec38",
  1667 => x"8156b497",
  1668 => x"04ff1454",
  1669 => x"73c83881",
  1670 => x"ff0bd40c",
  1671 => x"81ff0bd4",
  1672 => x"0cd00870",
  1673 => x"8f2a7081",
  1674 => x"06515153",
  1675 => x"72f33872",
  1676 => x"d00c7580",
  1677 => x"d3980c02",
  1678 => x"98050d04",
  1679 => x"02e8050d",
  1680 => x"77797b58",
  1681 => x"55558053",
  1682 => x"727625a3",
  1683 => x"38747081",
  1684 => x"055680f5",
  1685 => x"2d747081",
  1686 => x"055680f5",
  1687 => x"2d525271",
  1688 => x"712e8638",
  1689 => x"8151b4f1",
  1690 => x"04811353",
  1691 => x"b4c80480",
  1692 => x"517080d3",
  1693 => x"980c0298",
  1694 => x"050d0402",
  1695 => x"ec050d76",
  1696 => x"5574802e",
  1697 => x"80c4389a",
  1698 => x"1580e02d",
  1699 => x"5180c39a",
  1700 => x"2d80d398",
  1701 => x"0880d398",
  1702 => x"0880dab8",
  1703 => x"0c80d398",
  1704 => x"08545480",
  1705 => x"da940880",
  1706 => x"2e9b3894",
  1707 => x"1580e02d",
  1708 => x"5180c39a",
  1709 => x"2d80d398",
  1710 => x"08902b83",
  1711 => x"fff00a06",
  1712 => x"70750751",
  1713 => x"537280da",
  1714 => x"b80c80da",
  1715 => x"b8085372",
  1716 => x"802e9d38",
  1717 => x"80da8c08",
  1718 => x"fe147129",
  1719 => x"80daa008",
  1720 => x"0580dabc",
  1721 => x"0c70842b",
  1722 => x"80da980c",
  1723 => x"54b69e04",
  1724 => x"80daa408",
  1725 => x"80dab80c",
  1726 => x"80daa808",
  1727 => x"80dabc0c",
  1728 => x"80da9408",
  1729 => x"802e8b38",
  1730 => x"80da8c08",
  1731 => x"842b53b6",
  1732 => x"990480da",
  1733 => x"ac08842b",
  1734 => x"537280da",
  1735 => x"980c0294",
  1736 => x"050d0402",
  1737 => x"d8050d80",
  1738 => x"0b80da94",
  1739 => x"0c8454b0",
  1740 => x"962d80d3",
  1741 => x"9808802e",
  1742 => x"973880d4",
  1743 => x"88528051",
  1744 => x"b3982d80",
  1745 => x"d3980880",
  1746 => x"2e8638fe",
  1747 => x"54b6d804",
  1748 => x"ff145473",
  1749 => x"8024d838",
  1750 => x"738d3880",
  1751 => x"cdc85186",
  1752 => x"c52d7355",
  1753 => x"bcae0480",
  1754 => x"56810b80",
  1755 => x"dac00c88",
  1756 => x"5380cddc",
  1757 => x"5280d4be",
  1758 => x"51b4bc2d",
  1759 => x"80d39808",
  1760 => x"762e0981",
  1761 => x"06893880",
  1762 => x"d3980880",
  1763 => x"dac00c88",
  1764 => x"5380cde8",
  1765 => x"5280d4da",
  1766 => x"51b4bc2d",
  1767 => x"80d39808",
  1768 => x"893880d3",
  1769 => x"980880da",
  1770 => x"c00c80da",
  1771 => x"c008802e",
  1772 => x"81823880",
  1773 => x"d7ce0b80",
  1774 => x"f52d80d7",
  1775 => x"cf0b80f5",
  1776 => x"2d71982b",
  1777 => x"71902b07",
  1778 => x"80d7d00b",
  1779 => x"80f52d70",
  1780 => x"882b7207",
  1781 => x"80d7d10b",
  1782 => x"80f52d71",
  1783 => x"0780d886",
  1784 => x"0b80f52d",
  1785 => x"80d8870b",
  1786 => x"80f52d71",
  1787 => x"882b0753",
  1788 => x"5f54525a",
  1789 => x"56575573",
  1790 => x"81abaa2e",
  1791 => x"0981068f",
  1792 => x"38755180",
  1793 => x"c2e92d80",
  1794 => x"d3980856",
  1795 => x"b89d0473",
  1796 => x"82d4d52e",
  1797 => x"883880cd",
  1798 => x"f451b8e9",
  1799 => x"0480d488",
  1800 => x"527551b3",
  1801 => x"982d80d3",
  1802 => x"98085580",
  1803 => x"d3980880",
  1804 => x"2e83fb38",
  1805 => x"885380cd",
  1806 => x"e85280d4",
  1807 => x"da51b4bc",
  1808 => x"2d80d398",
  1809 => x"088a3881",
  1810 => x"0b80da94",
  1811 => x"0cb8ef04",
  1812 => x"885380cd",
  1813 => x"dc5280d4",
  1814 => x"be51b4bc",
  1815 => x"2d80d398",
  1816 => x"08802e8b",
  1817 => x"3880ce88",
  1818 => x"5186c52d",
  1819 => x"b9ce0480",
  1820 => x"d8860b80",
  1821 => x"f52d5473",
  1822 => x"80d52e09",
  1823 => x"810680ce",
  1824 => x"3880d887",
  1825 => x"0b80f52d",
  1826 => x"547381aa",
  1827 => x"2e098106",
  1828 => x"bd38800b",
  1829 => x"80d4880b",
  1830 => x"80f52d56",
  1831 => x"547481e9",
  1832 => x"2e833881",
  1833 => x"547481eb",
  1834 => x"2e8c3880",
  1835 => x"5573752e",
  1836 => x"09810682",
  1837 => x"f93880d4",
  1838 => x"930b80f5",
  1839 => x"2d55748e",
  1840 => x"3880d494",
  1841 => x"0b80f52d",
  1842 => x"5473822e",
  1843 => x"86388055",
  1844 => x"bcae0480",
  1845 => x"d4950b80",
  1846 => x"f52d7080",
  1847 => x"da8c0cff",
  1848 => x"0580da90",
  1849 => x"0c80d496",
  1850 => x"0b80f52d",
  1851 => x"80d4970b",
  1852 => x"80f52d58",
  1853 => x"76057782",
  1854 => x"80290570",
  1855 => x"80da9c0c",
  1856 => x"80d4980b",
  1857 => x"80f52d70",
  1858 => x"80dab00c",
  1859 => x"80da9408",
  1860 => x"59575876",
  1861 => x"802e81b7",
  1862 => x"38885380",
  1863 => x"cde85280",
  1864 => x"d4da51b4",
  1865 => x"bc2d80d3",
  1866 => x"98088282",
  1867 => x"3880da8c",
  1868 => x"0870842b",
  1869 => x"80da980c",
  1870 => x"7080daac",
  1871 => x"0c80d4ad",
  1872 => x"0b80f52d",
  1873 => x"80d4ac0b",
  1874 => x"80f52d71",
  1875 => x"82802905",
  1876 => x"80d4ae0b",
  1877 => x"80f52d70",
  1878 => x"84808029",
  1879 => x"1280d4af",
  1880 => x"0b80f52d",
  1881 => x"7081800a",
  1882 => x"29127080",
  1883 => x"dab40c80",
  1884 => x"dab00871",
  1885 => x"2980da9c",
  1886 => x"08057080",
  1887 => x"daa00c80",
  1888 => x"d4b50b80",
  1889 => x"f52d80d4",
  1890 => x"b40b80f5",
  1891 => x"2d718280",
  1892 => x"290580d4",
  1893 => x"b60b80f5",
  1894 => x"2d708480",
  1895 => x"80291280",
  1896 => x"d4b70b80",
  1897 => x"f52d7098",
  1898 => x"2b81f00a",
  1899 => x"06720570",
  1900 => x"80daa40c",
  1901 => x"fe117e29",
  1902 => x"770580da",
  1903 => x"a80c5259",
  1904 => x"5243545e",
  1905 => x"51525952",
  1906 => x"5d575957",
  1907 => x"bca70480",
  1908 => x"d49a0b80",
  1909 => x"f52d80d4",
  1910 => x"990b80f5",
  1911 => x"2d718280",
  1912 => x"29057080",
  1913 => x"da980c70",
  1914 => x"a02983ff",
  1915 => x"0570892a",
  1916 => x"7080daac",
  1917 => x"0c80d49f",
  1918 => x"0b80f52d",
  1919 => x"80d49e0b",
  1920 => x"80f52d71",
  1921 => x"82802905",
  1922 => x"7080dab4",
  1923 => x"0c7b7129",
  1924 => x"1e7080da",
  1925 => x"a80c7d80",
  1926 => x"daa40c73",
  1927 => x"0580daa0",
  1928 => x"0c555e51",
  1929 => x"51555580",
  1930 => x"51b4fb2d",
  1931 => x"81557480",
  1932 => x"d3980c02",
  1933 => x"a8050d04",
  1934 => x"02ec050d",
  1935 => x"7670872c",
  1936 => x"7180ff06",
  1937 => x"55565480",
  1938 => x"da94088a",
  1939 => x"3873882c",
  1940 => x"7481ff06",
  1941 => x"545580d4",
  1942 => x"885280da",
  1943 => x"9c081551",
  1944 => x"b3982d80",
  1945 => x"d3980854",
  1946 => x"80d39808",
  1947 => x"802eba38",
  1948 => x"80da9408",
  1949 => x"802e9b38",
  1950 => x"72842980",
  1951 => x"d4880570",
  1952 => x"08525380",
  1953 => x"c2e92d80",
  1954 => x"d39808f0",
  1955 => x"0a0653bd",
  1956 => x"a7047210",
  1957 => x"80d48805",
  1958 => x"7080e02d",
  1959 => x"525380c3",
  1960 => x"9a2d80d3",
  1961 => x"98085372",
  1962 => x"547380d3",
  1963 => x"980c0294",
  1964 => x"050d0402",
  1965 => x"e0050d79",
  1966 => x"70842c80",
  1967 => x"dabc0805",
  1968 => x"718f0652",
  1969 => x"5553728a",
  1970 => x"3880d488",
  1971 => x"527351b3",
  1972 => x"982d72a0",
  1973 => x"2980d488",
  1974 => x"05548074",
  1975 => x"80f52d56",
  1976 => x"5374732e",
  1977 => x"83388153",
  1978 => x"7481e52e",
  1979 => x"81f43881",
  1980 => x"70740654",
  1981 => x"5872802e",
  1982 => x"81e8388b",
  1983 => x"1480f52d",
  1984 => x"70832a79",
  1985 => x"06585676",
  1986 => x"9b3880d1",
  1987 => x"dc085372",
  1988 => x"89387280",
  1989 => x"d8880b81",
  1990 => x"b72d7680",
  1991 => x"d1dc0c73",
  1992 => x"53bfe404",
  1993 => x"758f2e09",
  1994 => x"810681b6",
  1995 => x"38749f06",
  1996 => x"8d2980d7",
  1997 => x"fb115153",
  1998 => x"811480f5",
  1999 => x"2d737081",
  2000 => x"055581b7",
  2001 => x"2d831480",
  2002 => x"f52d7370",
  2003 => x"81055581",
  2004 => x"b72d8514",
  2005 => x"80f52d73",
  2006 => x"70810555",
  2007 => x"81b72d87",
  2008 => x"1480f52d",
  2009 => x"73708105",
  2010 => x"5581b72d",
  2011 => x"891480f5",
  2012 => x"2d737081",
  2013 => x"055581b7",
  2014 => x"2d8e1480",
  2015 => x"f52d7370",
  2016 => x"81055581",
  2017 => x"b72d9014",
  2018 => x"80f52d73",
  2019 => x"70810555",
  2020 => x"81b72d92",
  2021 => x"1480f52d",
  2022 => x"73708105",
  2023 => x"5581b72d",
  2024 => x"941480f5",
  2025 => x"2d737081",
  2026 => x"055581b7",
  2027 => x"2d961480",
  2028 => x"f52d7370",
  2029 => x"81055581",
  2030 => x"b72d9814",
  2031 => x"80f52d73",
  2032 => x"70810555",
  2033 => x"81b72d9c",
  2034 => x"1480f52d",
  2035 => x"73708105",
  2036 => x"5581b72d",
  2037 => x"9e1480f5",
  2038 => x"2d7381b7",
  2039 => x"2d7780d1",
  2040 => x"dc0c8053",
  2041 => x"7280d398",
  2042 => x"0c02a005",
  2043 => x"0d0402cc",
  2044 => x"050d7e60",
  2045 => x"5e5a800b",
  2046 => x"80dab808",
  2047 => x"80dabc08",
  2048 => x"595c5680",
  2049 => x"5880da98",
  2050 => x"08782e81",
  2051 => x"bc38778f",
  2052 => x"06a01757",
  2053 => x"54739138",
  2054 => x"80d48852",
  2055 => x"76518117",
  2056 => x"57b3982d",
  2057 => x"80d48856",
  2058 => x"807680f5",
  2059 => x"2d565474",
  2060 => x"742e8338",
  2061 => x"81547481",
  2062 => x"e52e8181",
  2063 => x"38817075",
  2064 => x"06555c73",
  2065 => x"802e80f5",
  2066 => x"388b1680",
  2067 => x"f52d9806",
  2068 => x"597880e9",
  2069 => x"388b537c",
  2070 => x"527551b4",
  2071 => x"bc2d80d3",
  2072 => x"980880d9",
  2073 => x"389c1608",
  2074 => x"5180c2e9",
  2075 => x"2d80d398",
  2076 => x"08841b0c",
  2077 => x"9a1680e0",
  2078 => x"2d5180c3",
  2079 => x"9a2d80d3",
  2080 => x"980880d3",
  2081 => x"9808881c",
  2082 => x"0c80d398",
  2083 => x"08555580",
  2084 => x"da940880",
  2085 => x"2e9a3894",
  2086 => x"1680e02d",
  2087 => x"5180c39a",
  2088 => x"2d80d398",
  2089 => x"08902b83",
  2090 => x"fff00a06",
  2091 => x"70165154",
  2092 => x"73881b0c",
  2093 => x"787a0c7b",
  2094 => x"5480c286",
  2095 => x"04811858",
  2096 => x"80da9808",
  2097 => x"7826fec6",
  2098 => x"3880da94",
  2099 => x"08802eb4",
  2100 => x"387a51bc",
  2101 => x"b82d80d3",
  2102 => x"980880d3",
  2103 => x"980880ff",
  2104 => x"fffff806",
  2105 => x"555b7380",
  2106 => x"fffffff8",
  2107 => x"2e963880",
  2108 => x"d39808fe",
  2109 => x"0580da8c",
  2110 => x"082980da",
  2111 => x"a0080557",
  2112 => x"80c08304",
  2113 => x"80547380",
  2114 => x"d3980c02",
  2115 => x"b4050d04",
  2116 => x"02f4050d",
  2117 => x"74700881",
  2118 => x"05710c70",
  2119 => x"0880da90",
  2120 => x"08065353",
  2121 => x"718f3888",
  2122 => x"130851bc",
  2123 => x"b82d80d3",
  2124 => x"98088814",
  2125 => x"0c810b80",
  2126 => x"d3980c02",
  2127 => x"8c050d04",
  2128 => x"02f0050d",
  2129 => x"75881108",
  2130 => x"fe0580da",
  2131 => x"8c082980",
  2132 => x"daa00811",
  2133 => x"720880da",
  2134 => x"90080605",
  2135 => x"79555354",
  2136 => x"54b3982d",
  2137 => x"0290050d",
  2138 => x"0402f405",
  2139 => x"0d747088",
  2140 => x"2a83fe80",
  2141 => x"06707298",
  2142 => x"2a077288",
  2143 => x"2b87fc80",
  2144 => x"80067398",
  2145 => x"2b81f00a",
  2146 => x"06717307",
  2147 => x"0780d398",
  2148 => x"0c565153",
  2149 => x"51028c05",
  2150 => x"0d0402f8",
  2151 => x"050d028e",
  2152 => x"0580f52d",
  2153 => x"74882b07",
  2154 => x"7083ffff",
  2155 => x"0680d398",
  2156 => x"0c510288",
  2157 => x"050d0402",
  2158 => x"f4050d74",
  2159 => x"76785354",
  2160 => x"52807125",
  2161 => x"97387270",
  2162 => x"81055480",
  2163 => x"f52d7270",
  2164 => x"81055481",
  2165 => x"b72dff11",
  2166 => x"5170eb38",
  2167 => x"807281b7",
  2168 => x"2d028c05",
  2169 => x"0d0402e8",
  2170 => x"050d7756",
  2171 => x"80705654",
  2172 => x"737624b6",
  2173 => x"3880da98",
  2174 => x"08742eae",
  2175 => x"387351bd",
  2176 => x"b32d80d3",
  2177 => x"980880d3",
  2178 => x"98080981",
  2179 => x"057080d3",
  2180 => x"9808079f",
  2181 => x"2a770581",
  2182 => x"17575753",
  2183 => x"53747624",
  2184 => x"893880da",
  2185 => x"98087426",
  2186 => x"d4387280",
  2187 => x"d3980c02",
  2188 => x"98050d04",
  2189 => x"02f0050d",
  2190 => x"80d39408",
  2191 => x"165180c3",
  2192 => x"e62d80d3",
  2193 => x"9808802e",
  2194 => x"a0388b53",
  2195 => x"80d39808",
  2196 => x"5280d888",
  2197 => x"5180c3b7",
  2198 => x"2d80dac4",
  2199 => x"08547380",
  2200 => x"2e873880",
  2201 => x"d8885173",
  2202 => x"2d029005",
  2203 => x"0d0402dc",
  2204 => x"050d8070",
  2205 => x"5a557480",
  2206 => x"d3940825",
  2207 => x"b43880da",
  2208 => x"9808752e",
  2209 => x"ac387851",
  2210 => x"bdb32d80",
  2211 => x"d3980809",
  2212 => x"81057080",
  2213 => x"d3980807",
  2214 => x"9f2a7605",
  2215 => x"811b5b56",
  2216 => x"547480d3",
  2217 => x"94082589",
  2218 => x"3880da98",
  2219 => x"087926d6",
  2220 => x"38805578",
  2221 => x"80da9808",
  2222 => x"2781e338",
  2223 => x"7851bdb3",
  2224 => x"2d80d398",
  2225 => x"08802e81",
  2226 => x"b43880d3",
  2227 => x"98088b05",
  2228 => x"80f52d70",
  2229 => x"842a7081",
  2230 => x"06771078",
  2231 => x"842b80d8",
  2232 => x"880b80f5",
  2233 => x"2d5c5c53",
  2234 => x"51555673",
  2235 => x"802e80ce",
  2236 => x"38741682",
  2237 => x"2b80c7c2",
  2238 => x"0b80d1e8",
  2239 => x"120c5477",
  2240 => x"75311080",
  2241 => x"dac81155",
  2242 => x"56907470",
  2243 => x"81055681",
  2244 => x"b72da074",
  2245 => x"81b72d76",
  2246 => x"81ff0681",
  2247 => x"16585473",
  2248 => x"802e8b38",
  2249 => x"9c5380d8",
  2250 => x"885280c6",
  2251 => x"b5048b53",
  2252 => x"80d39808",
  2253 => x"5280daca",
  2254 => x"165180c6",
  2255 => x"f3047416",
  2256 => x"822b80c4",
  2257 => x"b40b80d1",
  2258 => x"e8120c54",
  2259 => x"7681ff06",
  2260 => x"81165854",
  2261 => x"73802e8b",
  2262 => x"389c5380",
  2263 => x"d8885280",
  2264 => x"c6ea048b",
  2265 => x"5380d398",
  2266 => x"08527775",
  2267 => x"311080da",
  2268 => x"c8055176",
  2269 => x"5580c3b7",
  2270 => x"2d80c792",
  2271 => x"04749029",
  2272 => x"75317010",
  2273 => x"80dac805",
  2274 => x"515480d3",
  2275 => x"98087481",
  2276 => x"b72d8119",
  2277 => x"59748b24",
  2278 => x"a43880c5",
  2279 => x"b3047490",
  2280 => x"29753170",
  2281 => x"1080dac8",
  2282 => x"058c7731",
  2283 => x"57515480",
  2284 => x"7481b72d",
  2285 => x"9e14ff16",
  2286 => x"565474f3",
  2287 => x"3802a405",
  2288 => x"0d0402fc",
  2289 => x"050d80d3",
  2290 => x"94081351",
  2291 => x"80c3e62d",
  2292 => x"80d39808",
  2293 => x"802e8938",
  2294 => x"80d39808",
  2295 => x"51b4fb2d",
  2296 => x"800b80d3",
  2297 => x"940c80c4",
  2298 => x"ee2d9feb",
  2299 => x"2d028405",
  2300 => x"0d0402fc",
  2301 => x"050d7251",
  2302 => x"70fd2eb2",
  2303 => x"3870fd24",
  2304 => x"8b3870fc",
  2305 => x"2e80d038",
  2306 => x"80c8e104",
  2307 => x"70fe2eb9",
  2308 => x"3870ff2e",
  2309 => x"09810680",
  2310 => x"c83880d3",
  2311 => x"94085170",
  2312 => x"802ebe38",
  2313 => x"ff1180d3",
  2314 => x"940c80c8",
  2315 => x"e10480d3",
  2316 => x"9408f405",
  2317 => x"7080d394",
  2318 => x"0c517080",
  2319 => x"25a33880",
  2320 => x"0b80d394",
  2321 => x"0c80c8e1",
  2322 => x"0480d394",
  2323 => x"08810580",
  2324 => x"d3940c80",
  2325 => x"c8e10480",
  2326 => x"d394088c",
  2327 => x"0580d394",
  2328 => x"0c80c4ee",
  2329 => x"2d9feb2d",
  2330 => x"0284050d",
  2331 => x"0402fc05",
  2332 => x"0d800b80",
  2333 => x"d3940c80",
  2334 => x"c4ee2d9e",
  2335 => x"d92d80d3",
  2336 => x"980880d3",
  2337 => x"840c80d1",
  2338 => x"e051a191",
  2339 => x"2d028405",
  2340 => x"0d047180",
  2341 => x"dac40c04",
  2342 => x"00ffffff",
  2343 => x"ff00ffff",
  2344 => x"ffff00ff",
  2345 => x"ffffff00",
  2346 => x"4b455953",
  2347 => x"50312020",
  2348 => x"20202000",
  2349 => x"00000000",
  2350 => x"4b455953",
  2351 => x"50322020",
  2352 => x"20202000",
  2353 => x"00000000",
  2354 => x"3d3d2056",
  2355 => x"6964656f",
  2356 => x"70616320",
  2357 => x"666f7220",
  2358 => x"5a58444f",
  2359 => x"53203d3d",
  2360 => x"00000000",
  2361 => x"3d3d3d3d",
  2362 => x"3d3d3d3d",
  2363 => x"3d3d3d3d",
  2364 => x"3d3d3d3d",
  2365 => x"3d3d3d3d",
  2366 => x"3d3d3d3d",
  2367 => x"00000000",
  2368 => x"52657365",
  2369 => x"74000000",
  2370 => x"5363616e",
  2371 => x"6c696e65",
  2372 => x"73000000",
  2373 => x"53776170",
  2374 => x"206a6f79",
  2375 => x"73746963",
  2376 => x"6b730000",
  2377 => x"4c6f6164",
  2378 => x"20524f4d",
  2379 => x"20100000",
  2380 => x"45786974",
  2381 => x"00000000",
  2382 => x"436f6c6f",
  2383 => x"72206d6f",
  2384 => x"64653a20",
  2385 => x"436f6c6f",
  2386 => x"72000000",
  2387 => x"436f6c6f",
  2388 => x"72206d6f",
  2389 => x"64653a20",
  2390 => x"4d6f6e6f",
  2391 => x"6368726f",
  2392 => x"6d650000",
  2393 => x"436f6c6f",
  2394 => x"72206d6f",
  2395 => x"64653a20",
  2396 => x"47726565",
  2397 => x"6e207068",
  2398 => x"6f737068",
  2399 => x"6f720000",
  2400 => x"436f6c6f",
  2401 => x"72206d6f",
  2402 => x"64653a20",
  2403 => x"416d6265",
  2404 => x"72206d6f",
  2405 => x"6e6f6368",
  2406 => x"726f6d65",
  2407 => x"00000000",
  2408 => x"4d6f6465",
  2409 => x"3a204f64",
  2410 => x"79737365",
  2411 => x"79322028",
  2412 => x"4e545343",
  2413 => x"29000000",
  2414 => x"4d6f6465",
  2415 => x"3a205669",
  2416 => x"64656f70",
  2417 => x"61632028",
  2418 => x"50414c29",
  2419 => x"00000000",
  2420 => x"3d3d2056",
  2421 => x"6964656f",
  2422 => x"70616320",
  2423 => x"666f7220",
  2424 => x"5a58554e",
  2425 => x"4f203d3d",
  2426 => x"00000000",
  2427 => x"5a58554e",
  2428 => x"4f3a2073",
  2429 => x"696e676c",
  2430 => x"65206a6f",
  2431 => x"79737469",
  2432 => x"636b0000",
  2433 => x"5a58554e",
  2434 => x"4f3a2032",
  2435 => x"206a6f79",
  2436 => x"73746963",
  2437 => x"6b207370",
  2438 => x"6c697474",
  2439 => x"65720000",
  2440 => x"5a58554e",
  2441 => x"4f3a2032",
  2442 => x"206a6f79",
  2443 => x"73746963",
  2444 => x"6b205647",
  2445 => x"41324d00",
  2446 => x"524f4d20",
  2447 => x"6c6f6164",
  2448 => x"696e6720",
  2449 => x"6661696c",
  2450 => x"65640000",
  2451 => x"4f4b0000",
  2452 => x"496e6974",
  2453 => x"69616c69",
  2454 => x"7a696e67",
  2455 => x"20534420",
  2456 => x"63617264",
  2457 => x"0a000000",
  2458 => x"16200000",
  2459 => x"14200000",
  2460 => x"15200000",
  2461 => x"53442069",
  2462 => x"6e69742e",
  2463 => x"2e2e0a00",
  2464 => x"53442063",
  2465 => x"61726420",
  2466 => x"72657365",
  2467 => x"74206661",
  2468 => x"696c6564",
  2469 => x"210a0000",
  2470 => x"53444843",
  2471 => x"20657272",
  2472 => x"6f72210a",
  2473 => x"00000000",
  2474 => x"57726974",
  2475 => x"65206661",
  2476 => x"696c6564",
  2477 => x"0a000000",
  2478 => x"52656164",
  2479 => x"20666169",
  2480 => x"6c65640a",
  2481 => x"00000000",
  2482 => x"43617264",
  2483 => x"20696e69",
  2484 => x"74206661",
  2485 => x"696c6564",
  2486 => x"0a000000",
  2487 => x"46415431",
  2488 => x"36202020",
  2489 => x"00000000",
  2490 => x"46415433",
  2491 => x"32202020",
  2492 => x"00000000",
  2493 => x"4e6f2070",
  2494 => x"61727469",
  2495 => x"74696f6e",
  2496 => x"20736967",
  2497 => x"0a000000",
  2498 => x"42616420",
  2499 => x"70617274",
  2500 => x"0a000000",
  2501 => x"4261636b",
  2502 => x"00000000",
  2503 => x"00000002",
  2504 => x"00000002",
  2505 => x"000024c8",
  2506 => x"00000a54",
  2507 => x"00000002",
  2508 => x"000024e4",
  2509 => x"00000a54",
  2510 => x"00000002",
  2511 => x"00002500",
  2512 => x"0000037f",
  2513 => x"00000001",
  2514 => x"00002508",
  2515 => x"00000000",
  2516 => x"00000001",
  2517 => x"00002514",
  2518 => x"00000001",
  2519 => x"00000002",
  2520 => x"00002524",
  2521 => x"0000246d",
  2522 => x"00000003",
  2523 => x"000027a8",
  2524 => x"00000002",
  2525 => x"00000003",
  2526 => x"00002798",
  2527 => x"00000004",
  2528 => x"00000002",
  2529 => x"00002530",
  2530 => x"00000f76",
  2531 => x"00000000",
  2532 => x"00000000",
  2533 => x"00000000",
  2534 => x"00002538",
  2535 => x"0000254c",
  2536 => x"00002564",
  2537 => x"00002580",
  2538 => x"000025a0",
  2539 => x"000025b8",
  2540 => x"00000002",
  2541 => x"000025d0",
  2542 => x"00000a54",
  2543 => x"00000002",
  2544 => x"000024e4",
  2545 => x"00000a54",
  2546 => x"00000002",
  2547 => x"00002500",
  2548 => x"0000037f",
  2549 => x"00000001",
  2550 => x"00002508",
  2551 => x"00000000",
  2552 => x"00000001",
  2553 => x"00002514",
  2554 => x"00000001",
  2555 => x"00000002",
  2556 => x"00002524",
  2557 => x"0000246d",
  2558 => x"00000003",
  2559 => x"000027a8",
  2560 => x"00000002",
  2561 => x"00000003",
  2562 => x"00002798",
  2563 => x"00000004",
  2564 => x"00000003",
  2565 => x"00002834",
  2566 => x"00000003",
  2567 => x"00000002",
  2568 => x"00002530",
  2569 => x"00000f76",
  2570 => x"00000000",
  2571 => x"00000000",
  2572 => x"00000000",
  2573 => x"000025ec",
  2574 => x"00002604",
  2575 => x"00002620",
  2576 => x"00000004",
  2577 => x"00002638",
  2578 => x"00002840",
  2579 => x"00000004",
  2580 => x"0000264c",
  2581 => x"00002720",
  2582 => x"00000000",
  2583 => x"00000000",
  2584 => x"00000000",
  2585 => x"00000000",
  2586 => x"00000000",
  2587 => x"00000000",
  2588 => x"00000000",
  2589 => x"00000000",
  2590 => x"00000000",
  2591 => x"00000000",
  2592 => x"00000000",
  2593 => x"00000000",
  2594 => x"00000000",
  2595 => x"00000000",
  2596 => x"00000000",
  2597 => x"00000000",
  2598 => x"00000000",
  2599 => x"00000000",
  2600 => x"00000000",
  2601 => x"00000000",
  2602 => x"00000000",
  2603 => x"00000006",
  2604 => x"00000043",
  2605 => x"00000042",
  2606 => x"0000003b",
  2607 => x"0000004b",
  2608 => x"00000033",
  2609 => x"0000001d",
  2610 => x"0000001b",
  2611 => x"0000001c",
  2612 => x"00000023",
  2613 => x"0000002b",
  2614 => x"00000000",
  2615 => x"00000000",
  2616 => x"00000002",
  2617 => x"00002d48",
  2618 => x"00002234",
  2619 => x"00000002",
  2620 => x"00002d66",
  2621 => x"00002234",
  2622 => x"00000002",
  2623 => x"00002d84",
  2624 => x"00002234",
  2625 => x"00000002",
  2626 => x"00002da2",
  2627 => x"00002234",
  2628 => x"00000002",
  2629 => x"00002dc0",
  2630 => x"00002234",
  2631 => x"00000002",
  2632 => x"00002dde",
  2633 => x"00002234",
  2634 => x"00000002",
  2635 => x"00002dfc",
  2636 => x"00002234",
  2637 => x"00000002",
  2638 => x"00002e1a",
  2639 => x"00002234",
  2640 => x"00000002",
  2641 => x"00002e38",
  2642 => x"00002234",
  2643 => x"00000002",
  2644 => x"00002e56",
  2645 => x"00002234",
  2646 => x"00000002",
  2647 => x"00002e74",
  2648 => x"00002234",
  2649 => x"00000002",
  2650 => x"00002e92",
  2651 => x"00002234",
  2652 => x"00000002",
  2653 => x"00002eb0",
  2654 => x"00002234",
  2655 => x"00000004",
  2656 => x"00002714",
  2657 => x"00000000",
  2658 => x"00000000",
  2659 => x"00000000",
  2660 => x"000023f2",
  2661 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

