---------------------------------------------------------
--
-- PS2 Keycode look up table
-- converts 7 bit key code to ASCII
-- Address bit 7 = CAPS Lock
-- Address bit 8 = Shift
--
-- J.E.Kent
-- 18th Oct 2004
--
library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity key_slice is
    Port (
       addr : in  std_logic_vector (8 downto 0);
       data : out std_logic_vector (7 downto 0)
    );
end key_slice;

architecture key_rom of key_slice is
  constant width   : integer := 8;
  constant memsize : integer := 512;

  type rom_array is array(0 to memsize-1) of std_logic_vector(width-1 downto 0);

  constant rom_data : rom_array :=
  ( 
"00000000", --00
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001001",
"01100000",
"00000000", --0F
"00000000", --10
"00000000",
"00000000",
"00000000",
"00000000",
"01110001",
"00110001",
"00000000",
"00000000",
"00000000",
"01111010",
"01110011",
"01100001",
"01110111",
"00110010",
"00000000", --1F
"00000000", --20
"01100011",
"01111000",
"01100100",
"01100101",
"00110100",
"00110011",
"00000000",
"00000000",
"00100000",
"01110110",
"01100110",
"01110100",
"01110010",
"00110101",
"00000000", --2F
"00000000", --30
"01101110",
"01100010",
"01101000",
"01100111",
"01111001",
"00110110",
"00000000",
"00000000",
"00000000",
"01101101",
"01101010",
"01110101",
"00110111",
"00111000",
"00000000", --3F
"00000000", --40
"00101100",
"01101011",
"01101001",
"01101111",
"00110000",
"00111001",
"00000000",
"00000000",
"00101110",
"00101111", --4A - /
"01101100",
"00111011",
"01110000",
"00101101",
"00000000", --4F
"00000000", --50
"00000000",
"00100111",
"00000000",
"01011011",
"00111101", --55 - =
"00000000",
"00000000",
"00000000",
"00000000",
"00001101", --5A - Enter
"01011101",
"00000000",
"01011100",
"00000000",
"00000000", --5F
"00000000", --60
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001000", --66 - Backspace
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000", --6F
"00000000", --70
"01111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00011011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00101010",
"00000000",
"00000000",
"00000000", --7F
"00000000", --80
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001001",
"01111110",
"00000000",
"00000000", --90
"00000000",
"00000000",
"00000000",
"00000000",
"01010001",
"00110001",
"00000000",
"00000000",
"00000000",
"01011010",
"01010011",
"01000001",
"01010111",
"00110010",
"00000000",
"00000000", --A0
"01000011",
"01011000",
"01000100",
"01000101",
"00110100",
"00110011",
"00000000",
"00000000",
"00100000",
"01010110",
"01000110",
"01010100",
"01010010",
"00110101",
"00000000",
"00000000", --B0
"01001110",
"01000010",
"01001000",
"01000111",
"01011001",
"00110110",
"00000000",
"00000000",
"00000000",
"01001101",
"01001010",
"01010101",
"00110111",
"00111000",
"00000000",
"00000000", --C0
"00101100",
"01001011",
"01001001",
"01001111",
"00110000",
"00111001",
"00000000",
"00000000",
"00101110",
"00101111",
"01001100",
"00111011",
"01010000",
"00101101",
"00000000",
"00000000", --D0
"00000000",
"00100111",
"00000000",
"01011011",
"00111101",
"00000000",
"00000000",
"00000000",
"00000000",
"00001101",
"01011101",
"00000000",
"01011100",
"00000000",
"00000000",
"00000000", --E0
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000", --F0
"01111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00011011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000", --100
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001001",
"01111110",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01010001",
"00100001",
"00000000",
"00000000",
"00000000",
"01011010",
"01010011",
"01000001",
"01010111",
"01000000",
"00000000",
"00000000",
"01000011",
"01011000",
"01000100",
"01000101",
"00100100",
"00100011",
"00000000",
"00000000",
"00100000",
"01010110",
"01000110",
"01010100",
"01010010",
"00100101",
"00000000",
"00000000",
"01001110",
"01000010",
"01001000",
"01000111",
"01011001",
"01011110",
"00000000",
"00000000",
"00000000",
"01001101",
"01001010",
"01010101",
"00100110",
"00101010",
"00000000",
"00000000",
"00111100",
"01001011",
"01001001",
"01001111",
"00101001",
"00101000",
"00000000",
"00000000",
"00111110",
"00111111",
"01001100",
"00111010",
"01010000",
"01011111",
"00000000",
"00000000",
"00000000",
"00100010",
"00000000",
"01111011",
"00101011",
"00000000",
"00000000",
"00000000",
"00000000",
"00001101",
"01111101",
"00000000",
"01111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00011011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00101010",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001001",
"01100000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01110001",
"00100001",
"00000000",
"00000000",
"00000000",
"01111010",
"01110011",
"01100001",
"01110111",
"01000000",
"00000000",
"00000000",
"01100011",
"01111000",
"01100100",
"01100101",
"00100100",
"00100011",
"00000000",
"00000000",
"00100000",
"01110110",
"01100110",
"01110100",
"01110010",
"00100101",
"00000000",
"00000000",
"01101110",
"01100010",
"01101000",
"01100111",
"01111001",
"01011110",
"00000000",
"00000000",
"00000000",
"01101101",
"01101010",
"01110101",
"00100110",
"00101010",
"00000000",
"00000000",
"00111100",
"01101011",
"01101001",
"01101111",
"00101001",
"00101000",
"00000000",
"00000000",
"00111110",
"00111111",
"01101100",
"00111010",
"01110000",
"01011111",
"00000000",
"00000000",
"00000000",
"00100010",
"00000000",
"01111011",
"00101011",
"00000000",
"00000000",
"00000000",
"00000000",
"00001101",
"01111101",
"00000000",
"01111100",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00001000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"01111111",
"00000000",
"00000000",
"00000000",
"00000000",
"00011011",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000",
"00000000"
  );
begin
   data <= rom_data(to_integer(unsigned(addr)));
end key_rom;
